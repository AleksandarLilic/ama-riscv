
`include "ama_riscv_defines.svh"
`include "ama_riscv_tb_defines.svh"

module ama_riscv_core_view (
    // top level signals
    input logic clk,
    input logic rst,
    rv_if_dc.TX dmem_req,
    input logic inst_retired,
    // internal signals
    input stage_ctrl_t ctrl_dec_exe,
    input stage_ctrl_t ctrl_exe_mem,
    input stage_ctrl_t ctrl_mem_wbk,
    input stage_ctrl_t ctrl_wbk_ret,
    input decoder_t decoded_exe,
    input branch_t branch_resolution_mem,
    input arch_width_t csr_tohost,
    input logic dc_stalled
);

// struct for all signals that are being tracked to retirement
typedef struct {
    inst_width_t inst;
    arch_width_t pc;
    logic branch_inst;
    logic branch_taken;
    logic bp_hit;
    arch_width_t dmem_addr;
    logic [3:0] dmem_size;
} retired_t;

pipeline_if_typed #(.T(inst_shadow_t)) inst_shadow ();
inst_shadow_t inst_shadow_ret;
pipeline_if_s nop ();
pipeline_if_s flush ();
retired_t r;

function automatic inst_shadow_t classify_inst(input inst_width_t inst);
    inst_shadow_t d;
    // d = 0; // to avoid X in wave, but Xs are easier to visually separate imo
    unique case (get_opc7(inst))
        OPC7_R_TYPE: d.r_type = inst;
        OPC7_I_TYPE,
        OPC7_LOAD,
        OPC7_JALR,
        OPC7_SYSTEM: d.i_type = inst;
        OPC7_STORE: d.s_type = inst;
        OPC7_BRANCH: d.b_type = inst;
        OPC7_JAL: d.j_type = inst;
        OPC7_LUI,
        OPC7_AUIPC: d.u_type = inst;
        // default: d = 0; // would catch flush as 0s inst ...
        default: ; // ... but make it Xs
    endcase
    return d;
endfunction

always_comb begin
    inst_shadow.dec = classify_inst(inst.dec);
    inst_shadow.exe = classify_inst(inst.exe);
    inst_shadow.mem = classify_inst(inst.mem);
    inst_shadow.wbk = classify_inst(inst.wbk);
    inst_shadow_ret = classify_inst(inst.ret);

    nop.dec = (inst.dec == `NOP);
    nop.exe = (inst.exe == `NOP);
    nop.mem = (inst.mem == `NOP);
    nop.wbk = (inst.wbk == `NOP);

    flush.dec = (inst.dec == 'h0);
    flush.exe = (inst.exe == 'h0);
    flush.mem = (inst.mem == 'h0);
    flush.wbk = (inst.wbk == 'h0);
end

// signals for tracing

// inst, pc
assign r.inst = inst.ret & {INST_WIDTH{inst_retired}};
assign r.pc = pc.ret & {ARCH_WIDTH{inst_retired}};

// branches
logic branch_inst_mem, branch_inst_wbk;
`STAGE(ctrl_exe_mem, 1'b1, decoded_exe.itype.branch, branch_inst_mem, 'h0)
`STAGE(ctrl_mem_wbk, 1'b1, branch_inst_mem, branch_inst_wbk, 'h0)
`STAGE(ctrl_wbk_ret, 1'b1, branch_inst_wbk, r.branch_inst, 'h0)

logic branch_taken_mem, branch_taken_wbk;
assign branch_taken_mem = ((branch_resolution_mem == B_T) && branch_inst_mem);
`STAGE(ctrl_mem_wbk, 1'b1, branch_taken_mem, branch_taken_wbk, 'h0)
`STAGE(ctrl_wbk_ret, 1'b1, branch_taken_wbk, r.branch_taken, 'h0)

`ifdef USE_BP
logic bp_hit_mem, bp_hit_wbk;
assign bp_hit_mem = (branch_inst_mem && `FE_CTRL.bp_hit);
`STAGE(ctrl_mem_wbk, 1'b1, bp_hit_mem, bp_hit_wbk, 'h0)
`STAGE(ctrl_wbk_ret, 1'b1, bp_hit_wbk, r.bp_hit, 'h0)
`else
assign r.bp_hit = 1'b0; // just to make trace function happy
`endif

arch_width_t csr_tohost_mem, csr_tohost_wbk;
`DFF_CI_RI_RVI(csr_tohost, csr_tohost_mem)
`DFF_CI_RI_RVI(csr_tohost_mem, csr_tohost_wbk)

// dmem
arch_width_t dmem_addr_exe, dmem_addr_mem, dmem_addr_wbk;
assign dmem_addr_exe = dmem_req.addr & {ARCH_WIDTH{dmem_req.valid}};

// enum class dmem_size_t {
//     lb, lh, lw, ld,
//     sb, sh, sw, sd,
//     no_access
// };
localparam int unsigned DMEM_SIZE_NA = 8;
logic [2:0] dmem_size;
logic [3:0] dmem_size_exe, dmem_size_mem, dmem_size_wbk;
assign dmem_size = dmem_req.dtype | {dmem_req.rtype, 2'b00};
assign dmem_size_exe = dmem_req.valid ? {1'b0, dmem_size} : DMEM_SIZE_NA;

`STAGE(ctrl_exe_mem, 1'b1, dmem_addr_exe, dmem_addr_mem, 'h0)
`STAGE(ctrl_mem_wbk, 1'b1, dmem_addr_mem, dmem_addr_wbk, 'h0)
`STAGE(ctrl_wbk_ret, 1'b1, dmem_addr_wbk, r.dmem_addr, 'h0)

`STAGE(ctrl_exe_mem, 1'b1, dmem_size_exe, dmem_size_mem, 'h0)
`STAGE(ctrl_mem_wbk, 1'b1, dmem_size_mem, dmem_size_wbk, DMEM_SIZE_NA)
`STAGE(ctrl_wbk_ret, 1'b1, dmem_size_wbk, r.dmem_size, DMEM_SIZE_NA)

// track down bubble
pipeline_if_s bubble ();
`DFF_CI_RI_RVI_EN(ctrl_dec_exe.en, ctrl_dec_exe.bubble, bubble.exe);
`DFF_CI_RI_RVI_EN(
    ctrl_exe_mem.en,
    (ctrl_exe_mem.bubble || bubble.exe),
    bubble.mem
);
`DFF_CI_RI_RVI_EN(ctrl_mem_wbk.en,
    (ctrl_mem_wbk.bubble || bubble.mem),
    bubble.wbk
);

endmodule
